module alu
(
   	 input      [4:0] rs, rt, 
   	 input      [4:0] rd,
	 input	    [4:0] shamt, 
	 input	    [5:0] funct
);
wire [31:0]sub_r;
wire [31:0]srl_r;
wire [31:0]add_r;


srl u2(rt, shamt, srl_r);
add u0(rs, rt, add_r);
sub u1(rs, rt, sub_r);

mux u3(add_r, sub_r, srl_r, funct, rd);

endmodule